`define VGA_WIDTH 640
`define VGA_HEIGHT 480

`define TEMPLATE_WIDTH 3
`define BOX_WIDTH 10
`define SEARCH_WIDTH 100


`define WHITE 4'hf

