`define VGA_WIDTH 640
`define VGA_HEIGHT 480

`define TEMPLATE_WIDTH 24
`define BOX_WIDTH 16
`define SEARCH_WIDTH 50

`define WHITE 4'hf

`define MAX_THRESHOLD 50